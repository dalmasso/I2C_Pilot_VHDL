----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:06:33 01/28/2014 
-- Design Name: 
-- Module Name:    porte_et - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity porte_et is
    Port ( sig1 : in  STD_LOGIC;
           sig2 : in  STD_LOGIC;
           sig_out : out  STD_LOGIC);
end porte_et;

architecture Behavioral of porte_et is
begin

sig_out <= sig1 and sig2;
			  
end Behavioral;

